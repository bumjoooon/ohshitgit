module tb;

initial begin

end

endmodule
