module tb;

initial begin

    tetstsetsetse salfjlkasf;
end

endmodule
