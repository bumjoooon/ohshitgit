module tb;

initial begin

    int a;
    int b;
    int c;
    reg [7:0] q;

end

endmodule
