module tb;

initial begin

    int a;
    int b;
    int c;
end

endmodule
